LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL; 
ENTITY final IS
	PORT(
		CLOCK_50 	: IN STD_LOGIC; -- 50MHz
		KEY			: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		-- LCD controller stuff
      LCD_RS, LCD_EN         : OUT STD_LOGIC;
      LCD_RW                 : OUT STD_LOGIC;
      LCD_ON                 : OUT STD_LOGIC;
      LCD_DATA               : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END final;

ARCHITECTURE arch OF final IS
		
	-- LCD display controller
	COMPONENT LCD_Display IS
		PORT( 
		 KEY         : IN STD_LOGIC_VECTOR(0 downto 0);
       CLOCK_50       : IN  STD_LOGIC;
       LCD_RS, LCD_EN         : OUT STD_LOGIC;
       LCD_RW                 : OUT   STD_LOGIC;
       LCD_ON                 : OUT STD_LOGIC;
       LCD_DATA               : INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		 GAME0 						: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		 GAME1 						: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		 GAME2 						: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		 GAME3 						: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		 OFFSET						: IN INTEGER RANGE 0 TO 3);
	END COMPONENT;
	
	COMPONENT ARROW_GENERATOR IS

	PORT(
		CLOCK		: IN  STD_LOGIC;
		RESET 	: IN 	STD_LOGIC;
	 	GAME0 	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		GAME1 	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		GAME2 	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		GAME3 	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0));

	END COMPONENT;
	
	
	SIGNAL COUNTER : INTEGER RANGE 0 TO 20000000:= 0;
	SIGNAL COUNTER2 : INTEGER RANGE 0 TO 5000000:= 0;
	
	SIGNAL reset: STD_LOGIC; 
	SIGNAL A0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL A1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL A2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL A3 : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL CLOCK :STD_LOGIC;
	SIGNAL CLOCK2: STD_LOGIC;
	
	SIGNAL OFFSET : INTEGER RANGE 0 TO 3:= 0;
	
BEGIN
	reset <= NOT KEY(1);
	--CLOCK <= KEY(0);
	
	PROCESS (CLOCK_50) -- 2.5 Hz clock
	BEGIN
		IF (rising_edge(CLOCK_50)) THEN
			COUNTER <= COUNTER + 1;
			IF (COUNTER <= 10000000) THEN
				CLOCK <= '1';
			ELSE
				CLOCK <= '0';
			END IF;
			
		END IF;		
	END PROCESS;
	
	PROCESS (CLOCK_50) -- 10 Hz clock
	BEGIN
		IF (rising_edge(CLOCK_50)) THEN
			COUNTER2 <= COUNTER2 + 1;
			IF (COUNTER2 <= 2500000) THEN
				CLOCK2 <= '1';
			ELSE
				CLOCK2 <= '0';
			END IF;
			
		END IF;		
	END PROCESS;
	
	PROCESS (CLOCK2)
	BEGIN
		IF (rising_edge(CLOCK2)) THEN
			OFFSET <= OFFSET + 1;
		END IF;
	
	END PROCESS;
	
	-- instantiate LCD controller
	lcd : LCD_Display PORT MAP(KEY(0 DOWNTO 0),CLOCK_50,LCD_RS, LCD_EN,LCD_RW ,LCD_ON,LCD_DATA, A0, A1, A2, A3,OFFSET);
	
	AG : ARROW_GENERATOR PORT MAP(CLOCK, reset, A0, A1, A2, A3);
END arch;